`include "c432.v"
module top;
reg N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
wire N223,N329,N370,N421,N430,N431,N432;
c432 m0(N1,N4,N8,N11,N14,N17,N21,N24,N27,N30, N34,N37,N40,N43,N47,N50,N53,N56,N60,N63, N66,N69,N73,N76,N79,N82,N86,N89,N92,N95, N99,N102,N105,N108,N112,N115,N223,N329,N370,N421, N430,N431,N432);
initial begin
	N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b0 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b0 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b1 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b1 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b1 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b0 ; N108=1'b1 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b0 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b0 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b0 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b0 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b1 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b1 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b1 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b0 ; N102=1'b1 ; N105=1'b1 ; N108=1'b1 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b0 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b0 ; N108=1'b1 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b0 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b0 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b1 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b0 ; N105=1'b1 ; N108=1'b1 ; N112=1'b1 ; N115=1'b1 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b1 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b0 ; 
	#5 N1=1'b0 ; N4=1'b0 ; N8=1'b0 ; N11=1'b0 ; N14=1'b0 ; N17=1'b0 ; N21=1'b0 ; N24=1'b0 ; N27=1'b0 ; N30=1'b0 ; N34=1'b0 ; N37=1'b0 ; N40=1'b0 ; N43=1'b0 ; N47=1'b0 ; N50=1'b0 ; N53=1'b0 ; N56=1'b0 ; N60=1'b0 ; N63=1'b0 ; N66=1'b0 ; N69=1'b0 ; N73=1'b0 ; N76=1'b0 ; N79=1'b0 ; N82=1'b0 ; N86=1'b0 ; N89=1'b0 ; N92=1'b0 ; N95=1'b0 ; N99=1'b1 ; N102=1'b1 ; N105=1'b0 ; N108=1'b0 ; N112=1'b0 ; N115=1'b1 ; 
end

initial begin
$monitor ($time, ": N1=%b N4=%b N8=%b N11=%b N14=%b N17=%b N21=%b N24=%b N27=%b N30=%b              N34=%b N37=%b N40=%b N43=%b N47=%b N50=%b N53=%b N56=%b N60=%b N63=%b              N66=%b N69=%b N73=%b N76=%b N79=%b N82=%b N86=%b N89=%b N92=%b N95=%b              N99=%b N102=%b N105=%b N108=%b N112=%b N115=%b N223=%b N329=%b N370=%b N421=%b              N430=%b N431=%b N432=%b ",N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,             N430,N431,N432);
$dumpfile("c432.vcd");
$dumpvars;
end

endmodule